          when others =>
                    instrOutput <= X"0000_0000";
		end case;
	end if;
end process;
end architecture;
